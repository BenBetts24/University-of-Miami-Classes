CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 71 640 760
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
30 C:\Circuit Maker\CM60S\BOM.DAT
0 7
0 71 640 760
144179219 0
0
6 Title:
5 Name:
0
0
0
6
10 Capacitor~
219 203 100 0 2 5
0 4 3
0
0 0 848 0
8 0.00001F
-29 -18 27 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8953 0 0
0
0
7 Ground~
168 308 167 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 116 82 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
11 Signal Gen~
195 71 65 0 19 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 1083179008 1036831949
20
1 1000 4.5 0.1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
8 4.4/4.6V
-29 -30 27 -22
2 V1
-7 -40 7 -32
0
0
41 %D %1 %2 DC 0 SIN(4.5 100m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
9 Resistor~
219 308 110 0 3 5
0 2 3 -1
0
0 0 880 90
4 100k
7 1 35 9
2 R2
13 -9 27 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
9 Resistor~
219 203 60 0 2 5
0 4 3
0
0 0 880 0
4 7.5k
-13 -14 15 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
6
0 2 3 0 0 4096 0 0 1 3 0 3
237 60
237 100
212 100
0 1 4 0 0 4096 0 0 1 5 0 3
168 60
168 100
194 100
2 2 3 0 0 4224 0 6 5 0 0 3
221 60
308 60
308 92
1 1 2 0 0 4224 0 5 2 0 0 2
308 128
308 161
1 1 4 0 0 4224 0 4 6 0 0 2
102 60
185 60
2 1 2 0 0 0 0 4 3 0 0 3
102 70
116 70
116 76
0
0
2073 0 1
0
0
0
0 0 0
0
0 0 0
10 2 1 80000
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2688158 1079360 100 100 0 0
0 0 0 0
428 189 589 259
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
1
168 60
0 4 0 0 1	0 2 0 0
2949288 8550976 100 100 0 0
77 66 587 246
640 71 1280 416
587 66
77 66
587 162
587 218
0 0
0.005 0 4.28 4.09333 0.005 0.005
12409 0
4 0.0005 2
2
155 60
0 4 0 0 1	0 5 0 0
302 60
0 3 0 0 1	0 3 0 0
3277660 4421696 100 100 0 0
77 66 587 246
640 416 1279 759
92 66
77 66
587 246
587 246
0 0
1765.71 1 -1.5 -1.5 75280.1 75280.1
12385 0
2 10000 0.5
2
158 60
0 4 0 0 1	0 5 0 0
300 60
0 3 0 0 1	0 3 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
