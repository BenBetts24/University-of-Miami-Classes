CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 71 640 760
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
30 C:\Circuit Maker\CM60S\BOM.DAT
0 7
0 71 640 760
144179219 0
0
6 Title:
5 Name:
0
0
0
18
11 Signal Gen~
195 70 361 0 64 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 1083179008 1036831949
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -1447456674
20
1 1000 4.5 0.1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
8 4.4/4.6V
-29 -30 27 -22
2 V3
-7 -40 7 -32
0
0
41 %D %1 %2 DC 0 SIN(4.5 100m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
7 Ground~
168 115 378 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 307 463 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
10 Capacitor~
219 281 356 0 2 5
0 4 3
0
0 0 848 0
4 100F
-14 -18 14 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
11 Signal Gen~
195 71 220 0 64 64
0 8 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 1083179008 1036831949
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -1447456674
20
1 1000 4.5 0.1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
8 4.4/4.6V
-29 -30 27 -22
2 V2
-7 -40 7 -32
0
0
41 %D %1 %2 DC 0 SIN(4.5 100m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
7 Ground~
168 116 237 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 308 322 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
10 Capacitor~
219 282 215 0 2 5
0 7 6
0
0 0 848 0
2 1F
-7 -18 7 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
10 Capacitor~
219 282 60 0 2 5
0 10 9
0
0 0 848 0
12 0.000000001F
-42 -18 42 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3549 0 0
0
0
7 Ground~
168 308 167 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
7 Ground~
168 116 82 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
11 Signal Gen~
195 71 65 0 19 64
0 11 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 1083179008 1036831949
20
1 1000 4.5 0.1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
8 4.4/4.6V
-29 -30 27 -22
2 V1
-7 -40 7 -32
0
0
41 %D %1 %2 DC 0 SIN(4.5 100m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
9 Resistor~
219 202 356 0 2 5
0 5 4
0
0 0 880 0
4 7.5k
-13 -14 15 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 307 406 0 3 5
0 2 3 -1
0
0 0 880 90
4 100k
7 0 35 8
2 R5
12 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 203 215 0 2 5
0 8 7
0
0 0 880 0
4 7.5k
-13 -14 15 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 308 265 0 3 5
0 2 6 -1
0
0 0 880 90
4 100k
7 0 35 8
2 R3
12 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 308 110 0 3 5
0 2 9 -1
0
0 0 880 90
4 100k
7 0 35 8
2 R2
12 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 203 60 0 2 5
0 11 10
0
0 0 880 0
4 7.5k
-13 -14 15 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
15
2 2 3 0 0 8320 0 4 14 0 0 3
290 356
307 356
307 388
2 1 4 0 0 4224 0 13 4 0 0 4
220 356
280 356
280 356
272 356
1 1 2 0 0 4224 0 14 3 0 0 2
307 424
307 457
1 1 5 0 0 4224 0 1 13 0 0 2
101 356
184 356
2 1 2 0 0 0 0 1 2 0 0 3
101 366
115 366
115 372
2 2 6 0 0 8320 0 8 16 0 0 3
291 215
308 215
308 247
2 1 7 0 0 4224 0 15 8 0 0 4
221 215
281 215
281 215
273 215
1 1 2 0 0 0 0 16 7 0 0 2
308 283
308 316
1 1 8 0 0 4224 0 5 15 0 0 2
102 215
185 215
2 1 2 0 0 0 0 5 6 0 0 3
102 225
116 225
116 231
2 2 9 0 0 8320 0 9 17 0 0 3
291 60
308 60
308 92
2 1 10 0 0 4224 0 18 9 0 0 4
221 60
281 60
281 60
273 60
1 1 2 0 0 0 0 17 10 0 0 2
308 128
308 161
1 1 11 0 0 4224 0 12 18 0 0 2
102 60
185 60
2 1 2 0 0 0 0 12 11 0 0 3
102 70
116 70
116 76
0
0
2073 0 1
0
0
0
0 0 0
0
0 0 0
10 2 1 80000
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2426008 1079360 100 100 0 0
0 0 0 0
443 203 604 273
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
1
167 60
0 11 0 0 1	0 14 0 0
3080558 8550976 100 100 0 0
77 66 587 246
640 71 1280 416
587 66
77 66
587 163
587 219
0 0
0.005 0 1.59 -0.09 0.005 0.005
12409 0
4 0.0005 2
2
155 60
0 11 0 0 1	0 14 0 0
302 60
0 9 0 0 1	0 11 0 0
2491094 4421696 100 100 0 0
77 66 587 246
640 419 1279 759
409 66
77 66
587 197
587 201
0 0
39059.8 1 -269.474 -296.842 75280.1 75280.1
12385 0
2 10000 200
4
158 60
0 11 0 0 1	0 14 0 0
300 60
0 9 0 0 1	0 11 0 0
300 215
0 6 0 0 1	0 6 0 0
300 356
0 3 0 0 1	0 1 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
